`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 11/24/2016 11:39:08 PM
// Design Name:
// Module Name: flipflop
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module flipflop(input logic in,clk,random,
                output logic out  );
   always_ff@(posedge clk)
       begin
        if(random == 1'b1)
            out<=in;
       end

endmodule
